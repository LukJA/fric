`ifndef _COMMON_VH_
`define _COMMON_VH_

package common;
    typedef enum logic { POS, NEG } sign_t;
endpackage

`endif // _COMMON_VH_
