package common;
    typedef enum logic {POS, NEG  } sign_t;
endpackage
